`timescale 1ns/1ps
`define clk_period 20

module tb_fma_top;

    parameter                       BW_EXP              =   8           ;
    parameter                       BW_MAN              =   9           ;
    parameter                       BW_FP               =   17          ;
    parameter                       BW_INT              =   8           ;
    parameter                       BW_ALIGN            =   9           ;
    parameter                       VALUE_MN            =   64          ;
    parameter                       M                   =   8           ;
    parameter                       N                   =   8           ;
    parameter                       K                   =   16          ;

    localparam                      HEAD_DIM            =   64          ;
    localparam                      HIDDEN_SIZE         =   2048        ;
    localparam                      INTERMEDIATE_SIZE   =   8192        ;

// instance signals
    reg                             clk                                 ;
    reg                             rst_n                               ;
    reg                             state_select                        ; //0:decode 1:prefill
    reg                             start_post_attn_norm_residual       ; //pulse,from PE
    reg                             start_post_attn_norm_sqrt           ; //pulse,from PE
    reg                             start1_norm1                        ;
    reg                             start1_sum_norm1                    ;
    reg                             start2_norm1                        ;
    reg                             start1_RoPE                         ;
    reg                             start2_RoPE                         ;
    reg     [VALUE_MN*BW_FP -1:0]   O_proj                              ; //8*4 pipeline,from PE
    reg     [VALUE_MN*BW_FP -1:0]   Z0                                  ; //8*4 from SRAM,512b
    reg     [VALUE_MN*BW_FP -1:0]   W_post_attn_norm                    ; //1*4 or 1*32 from SRAM,64*8b
    reg     [M*K*BW_FP      -1:0]   Input_norm1                         ; //8*16 ,from SRAM
    reg     [K*BW_FP        -1:0]   W_norm1                             ; //prefill 1*16     
    reg     [VALUE_MN*BW_FP -1:0]   QK_proj                             ; 
    reg     [VALUE_MN*BW_FP -1:0]   W_cos                               ; 
    reg     [VALUE_MN*BW_FP -1:0]   W_sin                               ; 
    reg     [VALUE_MN*BW_FP -1:0]   buffer_post_attn_norm_in            ; //from SRAM,512b
    wire    [M*K     *BW_FP   -1:0] buffer_norm1_out                    ; //to SRAM,512b
    wire    [VALUE_MN*2*BW_FP -1:0] buffer_post_attn_norm_out           ; //to SRAM,512b
    wire                            rms_result_valid                    ; // post_attn_norm
    wire                            scaled_x_valid                      ; // post_attn_norm
    wire    [VALUE_MN*2*BW_FP -1:0] buffer_RoPE                         ;
    wire                            busy_RoPE                           ;
    wire                            busy_post_attn_norm                 ;

    reg                             start_ffn_residual                  ;   // ffn_residual 
    reg       [VALUE_MN*BW_FP -1:0] D_proj                              ;   // ffn_residual 
    reg       [VALUE_MN*BW_FP -1:0] attn_residual_out                   ;   // ffn_residual
    wire                            busy_ffn_residual                   ;   // ffn_residual
    wire      [VALUE_MN*BW_FP -1:0] ffn_residual_out                    ;   // ffn_residual
    wire                            ffn_residual_out_valid              ;   // ffn_residual    

    reg                             start_ffn_mul                       ;   // ffn_mul
    reg       [VALUE_MN*BW_FP -1:0] U_proj                              ;   // ffn_mul
    reg       [VALUE_MN*BW_FP -1:0] silu_in                             ;   // ffn_mul
    wire                            busy_ffn_mul                        ;   // ffn_mul
    wire      [VALUE_MN*BW_FP -1:0] ffn_mul_out                         ;   // ffn_mul
    wire                            ffn_mul_out_valid                   ;   // ffn_mul

// general tb signals
    integer                         i,j                                 ;
    reg                             rope_start                          ;
    reg                             post_attn_norm_start                ;
    reg                             ffn_residual_start                  ;
    reg                             ffn_mul_start                       ;
    reg     [6:0]                   seq_len                             ;

// rope
    reg     [BW_FP - 1:0]           sin                     [0:4095]    ; 
    reg     [BW_FP - 1:0]           cos                     [0:4095]    ;
    reg     [BW_FP - 1:0]           k_origin                [0:4095]    ; 
    reg     [BW_FP - 1:0]           q_origin                [0:4095]    ;

    real                            q_FMA_dec               [0:4095]    ;
    real                            k_FMA_dec               [0:4095]    ; 

    reg     [2:0]                   rope_head_dim_cnt                   ;
    reg                             busy_RoPE_r                         ;
    wire                            busy_RoPE_fall                      ;
    reg                             RoPE_stage1                         ;
    reg                             RoPE_stage2                         ;
    reg                             RoPE_result_check                   ;

// post_attn_norm
    reg     [BW_FP - 1:0]           l0_input                [0:131071]  ; 
    reg     [BW_FP - 1:0]           l0_O_proj               [0:131071]  ;
    reg     [BW_FP - 1:0]           post_attn_norm_weight   [0:2047]    ; 

    reg                             busy_post_attn_norm_r               ;
    wire                            busy_post_attn_norm_fall            ;
    reg     [7:0]                   post_attn_norm_hidden_size_cnt      ;
    reg                             post_attn_norm_ready                ;
    reg     [BW_FP - 1:0]           scaled_x                [0:16383]   ; // 8 * 2048 = 16384
    reg     [3:0]                   post_attn_norm_seq_cnt              ; // seq 计数器  +1 表示 进8
    reg                             post_attn_norm_decode_flag          ;

    real                            post_attn_norm_result   [0:131071]  ; 

    real abs_error[0:63] ;
    real relative_error[0:63] ;
    real abs_error_temp;
    real relative_error_temp;

// ffn
// residual
    reg     [BW_FP - 1:0]           attn_residual_result        [0:131071]; 
    reg     [BW_FP - 1:0]           down_proj                   [0:131071];

    reg                             busy_ffn_residual_r                 ;
    wire                            busy_ffn_residual_fall              ;

    reg                             ffn_residual_ready                  ;
    reg     [7:0]                   ffn_residual_hidden_size_cnt        ;
    real                            ffn_residual_result   [0:131071]    ; // 8 * 2048 = 16384

    reg     [BW_FP - 1:0]           up_proj                     [0:524287];
    reg     [BW_FP - 1:0]           silu_gate                   [0:524287];

    reg                             busy_ffn_mul_r                 ;
    wire                            busy_ffn_mul_fall              ;

    reg                             ffn_mul_ready                  ;
    reg     [9:0]                   ffn_mul_intermediate_size_cnt  ;
    real                            ffn_mul_result   [0:524287]    ;

// FSM
    reg     [4:0]                   state, next_state                   ;
    // state
    localparam [4:0] 
        IDLE                            =   5'd0    ,
        ROPE_STAGE1                     =   5'd1    ,
        ROPE_STAGE2                     =   5'd2    ,
        ROPE_RESULT_SAVE                =   5'd3    ,
        POST_ATTN_NORM_RESIDUAL_PREFILL =   5'd4    ,
        POST_ATTN_NORM_SQRT             =   5'd5    ,
        POST_ATTN_NORM_PREFILL2DECODE   =   5'd6    ,
        POST_ATTN_NORM_RESIDUAL_DECODE  =   5'd7    ,
        POST_ATTN_NORM_RESULT_CHECK     =   5'd8    ,
        FFN_RESIDUAL                    =   5'd9    ,
        FFN_RESIDUAL_CHECK              =   5'd10   ,
        FFN_MUL                         =   5'd11   ,
        FFN_MUL_CHECK                   =   5'd12   ,
        STOP                            =   5'd31   ;

/******************** inst_fma_top *********************************/ 
    fma_top #(
        .BW_EXP  (BW_EXP  ),
        .BW_MAN  (BW_MAN  ),
        .BW_FP   (BW_FP   ),
        .BW_INT  (BW_INT  ),
        .BW_ALIGN(BW_ALIGN),
        .VALUE_MN(VALUE_MN),
        .M       (M       ),
        .N       (N       ),
        .K       (K       )
    )inst_fma_top(
        .clk                          (clk                          ),
        .rst_n                        (rst_n                        ),
        .state_select                 (state_select                 ),   //0:decode 1:prefill
        .start_post_attn_norm_residual(start_post_attn_norm_residual),   // post_attn_norm
        .start_post_attn_norm_sqrt    (start_post_attn_norm_sqrt    ),   // post_attn_norm
        .O_proj                       (O_proj                       ),   // post_attn_norm
        .Z0                           (Z0                           ),   // post_attn_norm
        .W_post_attn_norm             (W_post_attn_norm             ),   // post_attn_norm
        .buffer_post_attn_norm_in     (buffer_post_attn_norm_in     ),   // post_attn_norm
        .buffer_post_attn_norm_out    (buffer_post_attn_norm_out    ),   // post_attn_norm 
        .rms_result_valid             (rms_result_valid             ),   // post_attn_norm
        .scaled_x_valid               (scaled_x_valid               ),   // post_attn_norm
        .busy_post_attn_norm          (busy_post_attn_norm          ),   // post_attn_norm   
        .start1_norm1                 (start1_norm1                 ),
        .start1_sum_norm1             (start1_sum_norm1             ),
        .start2_norm1                 (start2_norm1                 ),
        .start1_RoPE                  (start1_RoPE                  ),   // RoPE
        .start2_RoPE                  (start2_RoPE                  ),   // RoPE
        .QK_proj                      (QK_proj                      ),   // RoPE 
        .W_cos                        (W_cos                        ),   // RoPE 
        .W_sin                        (W_sin                        ),   // RoPE 
        .buffer_RoPE                  (buffer_RoPE                  ),   // RoPE
        .busy_RoPE                    (busy_RoPE                    ),   // RoPE
        .Input_norm1                  (Input_norm1                  ),
        .W_norm1                      (W_norm1                      ),  
        .buffer_norm1_out             (buffer_norm1_out             ),
        .start_ffn_residual           (start_ffn_residual           ),   // ffn_residual 
        .D_proj                       (D_proj                       ),   // ffn_residual 
        .attn_residual_out            (attn_residual_out            ),   // ffn_residual
        .busy_ffn_residual            (busy_ffn_residual            ),   // ffn_residual
        .ffn_residual_out             (ffn_residual_out             ),   // ffn_residual
        .ffn_residual_out_valid       (ffn_residual_out_valid       ),   // ffn_residual    
        .start_ffn_mul                (start_ffn_mul                ),   // ffn_mul
        .U_proj                       (U_proj                       ),   // ffn_mul
        .silu_in                      (silu_in                      ),   // ffn_mul
        .busy_ffn_mul                 (busy_ffn_mul                 ),   // ffn_mul
        .ffn_mul_out                  (ffn_mul_out                  ),   // ffn_mul
        .ffn_mul_out_valid            (ffn_mul_out_valid            )    // ffn_mul
    );

/********************read and convert data*********************************/ 
    // rope
    // raw std BF16 storage
    reg [15:0]  sin_raw                     [0:4095]    ; 
    reg [15:0]  cos_raw                     [0:4095]    ;
    reg [15:0]  k_origin_raw                [0:4095]    ; 
    reg [15:0]  q_origin_raw                [0:4095]    ;
    reg [15:0]  k_rope_raw                  [0:4095]    ; 
    reg [15:0]  q_rope_raw                  [0:4095]    ;

    // std BF16 to Real storage
    real        sin_dec                     [0:4095]    ;
    real        cos_dec                     [0:4095]    ;
    real        k_origin_dec                [0:4095]    ;
    real        q_origin_dec                [0:4095]    ;
    real        k_rope_dec                  [0:4095]    ;
    real        q_rope_dec                  [0:4095]    ;

    // post_attn_norm
    reg [15:0]  l0_input_raw                [0:131071]  ;   // 64*2048=131072
    reg [15:0]  l0_O_proj_raw               [0:131071]  ;
    reg [15:0]  attn_residual_result_raw    [0:131071]  ; 
    reg [15:0]  post_attn_norm_result_raw   [0:131071]  ;
    reg [15:0]  post_attn_norm_weight_raw   [0:2047]    ; 

    // std BF16 to Real storage
    real        l0_input_dec                    [0:131071]  ;   // 64*2048=131072
    real        l0_O_proj_dec                   [0:131071]  ;
    real        attn_residual_result_dec        [0:131071]  ; 
    real        post_attn_norm_result_golden    [0:131071]  ;
    real        post_attn_norm_weight_dec       [0:2047]    ; 

    // ffn
    reg [15:0]  down_proj_raw                   [0:131071]  ;   // 64*2048=131072
    reg [15:0]  ffn_residual_result_raw         [0:131071]  ;
    reg [15:0]  up_proj_raw                     [0:524287]  ;   // 64*8192=524288
    reg [15:0]  silu_gate_raw                   [0:524287]  ;
    reg [15:0]  silu_dot_up_raw                 [0:524287]  ;

    real        down_proj_dec                   [0:131071]  ;
    real        ffn_residual_result_golden      [0:131071]  ;
    real        up_proj_dec                     [0:524287]  ;   // 64*8192=524288
    real        silu_golden                     [0:524287]  ;
    real        ffn_mul_golden                  [0:524287]  ;

    // $readmemb :loads a text file with binary values into a memory array
    initial begin
    // rope
        $readmemb("./rope_data/sin.txt", sin_raw);
        $readmemb("./rope_data/cos.txt", cos_raw);
        $readmemb("./rope_data/k_origin.txt", k_origin_raw);
        $readmemb("./rope_data/q_origin.txt", q_origin_raw);
        $readmemb("./rope_data/k_rope.txt", k_rope_raw);
        $readmemb("./rope_data/q_rope.txt", q_rope_raw);
    
    // post_attn_norm
        $readmemb("./layernorm_data/layer0_input_bf16.txt", l0_input_raw );
        $readmemb("./layernorm_data/layer0_attn_result_bf16.txt", l0_O_proj_raw );
        $readmemb("./layernorm_data/layer0_attn_residual_result_bf16.txt", attn_residual_result_raw);
        $readmemb("./layernorm_data/layer0_post_attention_layernorm_result_bf16.txt", post_attn_norm_result_raw );
        $readmemb("./layernorm_data/layer0_post_attention_layernorm_weight_bf16.txt", post_attn_norm_weight_raw );

    // ffn
        $readmemb("./ffn_data/down_proj_bf16.txt",down_proj_raw);
        $readmemb("./ffn_data/ffn_residual_result_bf16.txt",ffn_residual_result_raw);
        $readmemb("./ffn_data/up_proj_bf16.txt",up_proj_raw);
        $readmemb("./ffn_data/silu_gate_bf16.txt",silu_gate_raw);
        $readmemb("./ffn_data/silu_dot_up_bf16.txt",silu_dot_up_raw);


    // Convert std BF16 to Real
        for (i = 0; i < 4096; i = i + 1) begin
            sin_dec[i]      = std_bf16_to_dec(sin_raw[i]);
            cos_dec[i]      = std_bf16_to_dec(cos_raw[i]);
            k_origin_dec[i] = std_bf16_to_dec(k_origin_raw[i]);
            q_origin_dec[i] = std_bf16_to_dec(q_origin_raw[i]);
            k_rope_dec[i]   = std_bf16_to_dec(k_rope_raw[i]);
            q_rope_dec[i]   = std_bf16_to_dec(q_rope_raw[i]);
        end

        for (i = 0; i < 131072; i = i + 1) begin
            l0_input_dec[i]                 = std_bf16_to_dec(l0_input_raw[i]);
            l0_O_proj_dec[i]                = std_bf16_to_dec(l0_O_proj_raw[i]);
            attn_residual_result_dec[i]     = std_bf16_to_dec(attn_residual_result_raw[i]);
            post_attn_norm_result_golden[i] = std_bf16_to_dec(post_attn_norm_result_raw[i]);
            down_proj_dec[i]                = std_bf16_to_dec(down_proj_raw[i]);
            ffn_residual_result_golden[i]   = std_bf16_to_dec(ffn_residual_result_raw[i]);
        end

        for (i = 0; i < 2048; i = i + 1) begin
            post_attn_norm_weight_dec[i] = std_bf16_to_dec(post_attn_norm_weight_raw[i]);
        end

        for (i = 0; i < 524288; i = i + 1) begin
            up_proj_dec[i]       = std_bf16_to_dec(up_proj_raw[i]);
            silu_golden[i]       = std_bf16_to_dec(silu_gate_raw[i]);
            ffn_mul_golden[i]    = std_bf16_to_dec(silu_dot_up_raw[i]);
        end

        // Convert dec to BF16
        for (i = 0; i < 4096; i = i + 1) begin
            sin[i]      = dec_to_bf16(sin_dec[i]);
            cos[i]      = dec_to_bf16(cos_dec[i]);
            k_origin[i] = dec_to_bf16(k_origin_dec[i]);
            q_origin[i] = dec_to_bf16(q_origin_dec[i]);
        end

        for (i = 0; i < 131072; i = i + 1) begin
            l0_input[i]             = dec_to_bf16(l0_input_dec[i]);
            l0_O_proj[i]            = dec_to_bf16(l0_O_proj_dec[i]);
            attn_residual_result[i] = dec_to_bf16(attn_residual_result_dec[i]);
            down_proj[i]            = dec_to_bf16(down_proj_dec[i]);
        end

        for (i = 0; i < 2048; i = i + 1) begin
            post_attn_norm_weight[i] = dec_to_bf16(post_attn_norm_weight_dec[i]);
        end

        for (i = 0; i < 524288; i = i + 1) begin
            up_proj[i]     = dec_to_bf16(up_proj_dec[i]);
            silu_gate[i]   = dec_to_bf16(silu_golden[i]);
        end
    end

/******************** RoPE ****************************/ 
    // negedge edge detect
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) 
            busy_RoPE_r <= 1'b0;
        else 
            busy_RoPE_r <= busy_RoPE;
    end
    assign busy_RoPE_fall = busy_RoPE_r && !busy_RoPE;

/************************** post_attn_norm ****************************/ 
    // negedge edge detect
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) 
            busy_post_attn_norm_r <= 1'b0;
        else 
            busy_post_attn_norm_r <= busy_post_attn_norm;
    end
    assign busy_post_attn_norm_fall = busy_post_attn_norm_r && !busy_post_attn_norm;

    // 模拟sram 存储 rms 分子
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            for (i = 0; i < 16384; i = i + 1) begin
                scaled_x[i] <= 1'b0 ;
            end
        end
        else if (scaled_x_valid) begin
            if (state_select) begin
                for (i = 0; i < M; i = i + 1) begin
                    for (j = 0; j < N; j = j + 1) begin
                        scaled_x[HIDDEN_SIZE*i + j + post_attn_norm_hidden_size_cnt*N] <= buffer_post_attn_norm_out[N*(i+M)*BW_FP + j*BW_FP +: BW_FP] ;
                    end
                end
            end
            else begin
                if(!post_attn_norm_decode_flag) begin
                    for (j = 0; j < 64; j = j + 1) begin
                        scaled_x[j + post_attn_norm_hidden_size_cnt*64] <= buffer_post_attn_norm_out[(j+64)*BW_FP +: BW_FP] ;
                    end
                end 
            end
        end
    end

    // 模拟sram 存储 rms 结果
    always @(posedge clk or negedge rst_n) begin
        if (state_select) begin
            if (rms_result_valid & (post_attn_norm_seq_cnt > 0)) begin
                for (i = 0; i < M; i = i + 1) begin
                    for (j = 0; j < N; j = j + 1) begin
                        post_attn_norm_result[HIDDEN_SIZE*(i + (post_attn_norm_seq_cnt-1) * 8) + j + (post_attn_norm_hidden_size_cnt-1'd1)*N] = bf16_to_dec(buffer_post_attn_norm_out[N*i*BW_FP + j*BW_FP +: BW_FP]);
                        post_attn_norm_result[HIDDEN_SIZE*(i + (post_attn_norm_seq_cnt-1) * 8) + j + post_attn_norm_hidden_size_cnt*N] = bf16_to_dec(buffer_post_attn_norm_out[N*(i+M)*BW_FP + j*BW_FP +: BW_FP]);
                    end
                end
            end
        end
        else begin
            if(rms_result_valid & post_attn_norm_decode_flag) begin
                for (j = 0; j < 64; j = j + 1) begin
                    post_attn_norm_result[HIDDEN_SIZE*seq_len + j + (post_attn_norm_hidden_size_cnt-1'd1)*64] = bf16_to_dec(buffer_post_attn_norm_out[j*BW_FP +: BW_FP]);
                    post_attn_norm_result[HIDDEN_SIZE*seq_len + j + post_attn_norm_hidden_size_cnt*64] = bf16_to_dec(buffer_post_attn_norm_out[(j+64)*BW_FP +: BW_FP]);
                end
            end
        end
    end

/************************** ffn ****************************/ 
//ffn residual
    // negedge edge detect
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) 
            busy_ffn_residual_r <= 1'b0;
        else 
            busy_ffn_residual_r <= busy_ffn_residual;
    end
    assign busy_ffn_residual_fall = busy_ffn_residual_r && !busy_ffn_residual;

    // 模拟sram 存储 rms 结果
    always @(posedge clk or negedge rst_n) begin
        if (ffn_residual_out_valid) begin
            for (i = 0; i < M; i = i + 1) begin
                for (j = 0; j < N; j = j + 1) begin
                    ffn_residual_result[HIDDEN_SIZE*i + j + ffn_residual_hidden_size_cnt*N] = bf16_to_dec(ffn_residual_out[N*i*BW_FP + j*BW_FP +: BW_FP]);
                end
            end
        end
    end

//ffn mul
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) 
            busy_ffn_mul_r <= 1'b0;
        else 
            busy_ffn_mul_r <= busy_ffn_mul;
    end
    assign busy_ffn_mul_fall = busy_ffn_mul_r && !busy_ffn_mul;

    // 模拟sram 存储 rms 结果
    always @(posedge clk or negedge rst_n) begin
        if (ffn_mul_out_valid) begin
            for (i = 0; i < M; i = i + 1) begin
                for (j = 0; j < N; j = j + 1) begin
                    ffn_mul_result[INTERMEDIATE_SIZE*i + j + ffn_mul_intermediate_size_cnt*N] = bf16_to_dec(ffn_mul_out[N*i*BW_FP + j*BW_FP +: BW_FP]);
                end
            end
        end
    end
/******************** FSM ****************************/ 

    // update state
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) 
            state <= IDLE;
        else 
            state <= next_state;
    end

    // next state logic
    always @(*) begin
        case(state)
            IDLE: begin
                if(rope_start)
                    next_state = ROPE_STAGE1;
                else if(post_attn_norm_start)
                    next_state = POST_ATTN_NORM_RESIDUAL_PREFILL;
                else if(ffn_residual_start)
                    next_state = FFN_RESIDUAL;
                else if(ffn_mul_start)
                    next_state = FFN_MUL;
                else
                    next_state = IDLE;
            end
            ROPE_STAGE1:   
                next_state = busy_RoPE_fall ? ROPE_STAGE2 : ROPE_STAGE1 ;
            ROPE_STAGE2: 
                next_state = busy_RoPE_fall ? ROPE_RESULT_SAVE : ROPE_STAGE2 ;
            ROPE_RESULT_SAVE:
                next_state = STOP ;
            POST_ATTN_NORM_RESIDUAL_PREFILL : begin  
                if(busy_post_attn_norm_fall) begin
                    if(post_attn_norm_hidden_size_cnt == 8'd255)
                        next_state = POST_ATTN_NORM_SQRT ;
                    else
                        next_state = POST_ATTN_NORM_RESIDUAL_PREFILL ;
                end
                else
                    next_state = POST_ATTN_NORM_RESIDUAL_PREFILL ;
            end
            POST_ATTN_NORM_SQRT : begin
                if(busy_post_attn_norm_fall) begin
                    if(state_select) begin
                        if(post_attn_norm_seq_cnt * 8 >= seq_len)
                            next_state = POST_ATTN_NORM_PREFILL2DECODE ;
                        else
                            next_state = POST_ATTN_NORM_RESIDUAL_PREFILL ;
                    end
                    else
                        next_state = POST_ATTN_NORM_RESIDUAL_DECODE ;
                end
                else
                    next_state = POST_ATTN_NORM_SQRT;
            end
            POST_ATTN_NORM_PREFILL2DECODE : begin
                if(busy_post_attn_norm_fall) begin
                    if(post_attn_norm_hidden_size_cnt == 8'd255)
                        next_state = POST_ATTN_NORM_RESIDUAL_DECODE ;
                    else
                        next_state = POST_ATTN_NORM_PREFILL2DECODE ;
                end
                else
                    next_state = POST_ATTN_NORM_PREFILL2DECODE ;
            end
            POST_ATTN_NORM_RESIDUAL_DECODE : begin
                if(busy_post_attn_norm_fall) begin
                    if(post_attn_norm_hidden_size_cnt == 8'd31) begin
                        if(!post_attn_norm_decode_flag)
                            next_state = POST_ATTN_NORM_SQRT ;
                        else
                            next_state = POST_ATTN_NORM_RESULT_CHECK ;
                    end
                    else
                        next_state = POST_ATTN_NORM_RESIDUAL_DECODE ;
                end
                else
                    next_state = POST_ATTN_NORM_RESIDUAL_DECODE ;
            end
            POST_ATTN_NORM_RESULT_CHECK : next_state = STOP ;
            FFN_RESIDUAL : begin
                if(busy_ffn_residual_fall) begin
                    if(ffn_residual_hidden_size_cnt == 8'd255)
                        next_state = FFN_RESIDUAL_CHECK ;
                    else
                        next_state = FFN_RESIDUAL ;
                end
                else
                    next_state = FFN_RESIDUAL ;
            end
            FFN_RESIDUAL_CHECK : next_state = STOP ;
            FFN_MUL : begin
                if(busy_ffn_mul_fall) begin
                    if(ffn_mul_intermediate_size_cnt == 10'd1023)
                        next_state = FFN_MUL_CHECK ;
                    else
                        next_state = FFN_MUL ;
                end
                else
                    next_state = FFN_MUL ;
            end
            FFN_MUL_CHECK : next_state = STOP ;
            STOP:    next_state = IDLE;
            default: next_state = IDLE;
        endcase
    end

    // rope fsm control
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            // RoPE init
            start1_RoPE <= 1'b0;
            start2_RoPE <= 1'b0;
            QK_proj     <= 1'b0;
            W_cos       <= 1'b0;
            W_sin       <= 1'b0;
            rope_head_dim_cnt <= 1'b0;
            RoPE_stage1 <= 1'd0;
            RoPE_stage2 <= 1'd0;
        end 
        else begin
            case(state)
                IDLE: begin
                    // RoPE
                    start1_RoPE <= 1'b0;
                    start2_RoPE <= 1'b0;
                    QK_proj     <= 1'b0;
                    W_cos       <= 1'b0;
                    W_sin       <= 1'b0;
                    rope_head_dim_cnt <= 1'b0;
                    RoPE_stage1 <= 1'd0;
                    RoPE_stage2 <= 1'd0;
                end
            // RoPE
                ROPE_STAGE1 : begin
                    if(!RoPE_stage1) begin
                        RoPE_stage1 <= 1'b1;
                        RoPE_stage2 <= 1'b0;

                        start1_RoPE <= 1'b1;
                        for(i = 0; i < M ; i = i + 1) begin
                            for(j = 0; j < N; j = j + 1) begin
                                QK_proj[N*i*BW_FP + j*BW_FP +: BW_FP] <= q_origin[HEAD_DIM*i + j + rope_head_dim_cnt*N];
                                W_cos[N*i*BW_FP + j*BW_FP +: BW_FP]   <= cos[HEAD_DIM*i + j + rope_head_dim_cnt*N];
                                W_sin[N*i*BW_FP + j*BW_FP +: BW_FP]   <= sin[HEAD_DIM*i + j + rope_head_dim_cnt*N];
                            end
                        end
                    end
                    else begin
                        start1_RoPE <= 1'b0;
                    end
                end
                ROPE_STAGE2 : begin
                    if(!RoPE_stage2) begin
                        RoPE_stage1 <= 1'b0;
                        RoPE_stage2 <= 1'b1;

                        start2_RoPE <= 1'b1;
                        for(i = 0; i < M ; i = i + 1) begin
                            for(j = 0; j < N; j = j + 1) begin
                                QK_proj[N*i*BW_FP + j*BW_FP +: BW_FP] <= q_origin[HEAD_DIM*i + j + rope_head_dim_cnt*N + 4* N];
                                W_cos[N*i*BW_FP + j*BW_FP +: BW_FP]   <= cos[HEAD_DIM*i + j + rope_head_dim_cnt*N + 4* N];
                                W_sin[N*i*BW_FP + j*BW_FP +: BW_FP]   <= sin[HEAD_DIM*i + j + rope_head_dim_cnt*N + 4* N];
                            end
                        end
                    end
                    else begin
                        start2_RoPE <= 1'b0;
                    end
                end
                ROPE_RESULT_SAVE: begin
                    for(i = 0; i < M ; i = i + 1) begin
                        for(j = 0; j < N; j = j + 1) begin
                            q_FMA_dec[HEAD_DIM*i + j + rope_head_dim_cnt*N] = bf16_to_dec(buffer_RoPE[N*i*BW_FP + j*BW_FP +: BW_FP]);
                            $display("q_FMA_dec[%0d]: %f", HEAD_DIM*i + j + rope_head_dim_cnt*N, q_FMA_dec[HEAD_DIM*i + j + rope_head_dim_cnt*N]);
                            $display("q_rope_dec[%0d]: %f", HEAD_DIM*i + j + rope_head_dim_cnt*N, q_rope_dec[HEAD_DIM*i + j + rope_head_dim_cnt*N]);
                            q_FMA_dec[HEAD_DIM*i + j + rope_head_dim_cnt*N + 4* N] = bf16_to_dec(buffer_RoPE[N*(i+M)*BW_FP + j*BW_FP +: BW_FP]);
                        end
                    end
                end
                default : begin
                    // RoPE
                    start1_RoPE <= 1'b0;
                    start2_RoPE <= 1'b0;
                    QK_proj     <= 1'b0;
                    W_cos       <= 1'b0;
                    W_sin       <= 1'b0;
                    rope_head_dim_cnt <= 1'b0;
                    RoPE_stage1 <= 1'd0;
                    RoPE_stage2 <= 1'd0;
                    RoPE_result_check <= 1'd0;
                end
            endcase
        end
    end

    // post_attn_norm fsm control
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            seq_len <= 7'd16;
            post_attn_norm_hidden_size_cnt <= 1'b0;
            start_post_attn_norm_residual <= 1'b0;
            start_post_attn_norm_sqrt <= 1'b0;
            post_attn_norm_ready <= 1'b0;
            O_proj <= 1'b0;
            Z0 <= 1'b0;
            buffer_post_attn_norm_in <= 1'b0;
            W_post_attn_norm <= 1'b0;
            post_attn_norm_seq_cnt <= 1'b0;
            state_select <= 1'b1;
            post_attn_norm_decode_flag <= 1'b0;
        end 
        else begin
            case(state)
                IDLE: begin
                    seq_len <= 7'd16;
                    post_attn_norm_hidden_size_cnt <= 1'b0;
                    start_post_attn_norm_residual <= 1'b0;
                    start_post_attn_norm_sqrt <= 1'b0;
                    post_attn_norm_ready <= 1'b0;
                    O_proj <= 1'b0;
                    Z0 <= 1'b0;
                    buffer_post_attn_norm_in <= 1'b0;
                    W_post_attn_norm <= 1'b0;
                    post_attn_norm_seq_cnt <= 1'b0;
                    state_select <= 1'b1;
                    post_attn_norm_decode_flag <= 1'b0;
                end
                POST_ATTN_NORM_RESIDUAL_PREFILL : begin
                    if(!post_attn_norm_ready) begin
                        start_post_attn_norm_residual <= 1'b1;
                        post_attn_norm_ready <= 1'b1;
                        for(i = 0; i < M ; i = i + 1) begin
                            for(j = 0; j < N; j = j + 1) begin
                                O_proj[N*i*BW_FP + j*BW_FP +: BW_FP] <= l0_O_proj[HIDDEN_SIZE*(i + post_attn_norm_seq_cnt * 8) + j + post_attn_norm_hidden_size_cnt*N];
                                Z0[N*i*BW_FP + j*BW_FP +: BW_FP] <= l0_input[HIDDEN_SIZE*(i + post_attn_norm_seq_cnt * 8) + j + post_attn_norm_hidden_size_cnt*N];
                            end
                        end
                        for(j = 0; j < N; j = j + 1) begin
                            W_post_attn_norm[j*BW_FP +: BW_FP] <= post_attn_norm_weight[j + post_attn_norm_hidden_size_cnt*N];
                        end
                        if(post_attn_norm_seq_cnt == 8'd0) begin
                            for(i = 0; i < M ; i = i + 1) begin
                                for(j = 0; j < N; j = j + 1) begin
                                    buffer_post_attn_norm_in[N*i*BW_FP + j*BW_FP +: BW_FP] <= 1'b0;
                                end
                            end
                        end
                        else begin
                            for(i = 0; i < M ; i = i + 1) begin
                                for(j = 0; j < N; j = j + 1) begin
                                    buffer_post_attn_norm_in[N*i*BW_FP + j*BW_FP +: BW_FP] <= scaled_x[HIDDEN_SIZE*i+ j + post_attn_norm_hidden_size_cnt*N];
                                end
                            end
                        end
                    end
                    else if(busy_post_attn_norm_fall) begin
                        post_attn_norm_ready <= 1'd0;
                        post_attn_norm_hidden_size_cnt <= post_attn_norm_hidden_size_cnt + 1'd1;
                        if(post_attn_norm_hidden_size_cnt == 8'd255) begin
                            post_attn_norm_seq_cnt <= post_attn_norm_seq_cnt + 1'd1;
                        end
                    end
                    else begin
                        start_post_attn_norm_residual <= 1'b0;
                    end
                end
                POST_ATTN_NORM_SQRT: begin
                    if(!post_attn_norm_ready) begin
                        start_post_attn_norm_sqrt <= 1'b1;
                        post_attn_norm_ready <= 1'b1;
                    end
                    else if(busy_post_attn_norm_fall) begin
                        post_attn_norm_ready <= 1'd0;
                    end
                    else begin
                        start_post_attn_norm_sqrt <= 1'b0;
                    end
                end
                POST_ATTN_NORM_PREFILL2DECODE : begin
                    if(!post_attn_norm_ready) begin
                        start_post_attn_norm_residual <= 1'b1;
                        post_attn_norm_ready <= 1'b1;
                        O_proj <= 1'd0;
                        Z0 <= 1'd0;
                        W_post_attn_norm <= 1'd0;
                        for(i = 0; i < M ; i = i + 1) begin
                            for(j = 0; j < N; j = j + 1) begin
                                buffer_post_attn_norm_in[N*i*BW_FP + j*BW_FP +: BW_FP] <= scaled_x[HIDDEN_SIZE*i+ j + post_attn_norm_hidden_size_cnt*N];
                            end
                        end
                    end
                    else if(busy_post_attn_norm_fall) begin
                        post_attn_norm_ready <= 1'd0;
                        post_attn_norm_hidden_size_cnt <= post_attn_norm_hidden_size_cnt + 1'd1;
                        if(post_attn_norm_hidden_size_cnt == 8'd255) begin
                            state_select <= 1'd0;
                        end
                    end
                    else begin
                        start_post_attn_norm_residual <= 1'b0;
                    end
                end
                POST_ATTN_NORM_RESIDUAL_DECODE : begin
                    if(!post_attn_norm_ready) begin
                        start_post_attn_norm_residual <= 1'b1;
                        post_attn_norm_ready <= 1'b1;
                        if (!post_attn_norm_decode_flag) begin
                            for(j = 0; j < 64; j = j + 1) begin
                                O_proj[j*BW_FP +: BW_FP] <= l0_O_proj[HIDDEN_SIZE*seq_len + j + post_attn_norm_hidden_size_cnt*64];
                                Z0[j*BW_FP +: BW_FP] <= l0_input[HIDDEN_SIZE*seq_len+ j + post_attn_norm_hidden_size_cnt*64];
                                W_post_attn_norm[j*BW_FP +: BW_FP] <= post_attn_norm_weight[j + post_attn_norm_hidden_size_cnt*64];
                            end
                            buffer_post_attn_norm_in <= 1'b0;
                        end
                        else begin
                            O_proj <= 1'd0;
                            Z0 <= 1'd0;
                            W_post_attn_norm <= 1'd0;
                            for(j = 0; j < 64; j = j + 1) begin
                                buffer_post_attn_norm_in[j*BW_FP +: BW_FP] <= scaled_x[j + post_attn_norm_hidden_size_cnt*64];
                            end
                        end
                    end
                    else if(busy_post_attn_norm_fall) begin
                        post_attn_norm_ready <= 1'd0;
                        if(post_attn_norm_hidden_size_cnt >= 8'd31) begin
                            post_attn_norm_decode_flag <= ~post_attn_norm_decode_flag;
                            post_attn_norm_hidden_size_cnt <= 1'd0;
                            if(post_attn_norm_decode_flag)
                                seq_len <= seq_len + 1'd1;
                        end
                        else begin
                            post_attn_norm_hidden_size_cnt <= post_attn_norm_hidden_size_cnt + 1'd1;
                        end
                    end
                    else begin
                        start_post_attn_norm_residual <= 1'b0;
                    end
                end
                POST_ATTN_NORM_RESULT_CHECK: begin
                    for (i =0 ; i< seq_len; i = i + 1) begin
                        for(j = 0; j < 2048; j = j + 1) begin
                            $display("post_attn_norm_result_golden[%0d]: %f", i*2048+j, post_attn_norm_result_golden[i*2048+j]);
                            $display("post_attn_norm_result[%0d]: %f", i*2048+j, post_attn_norm_result[i*2048+j]);
                            abs_error_temp =abs_error_temp + $abs(post_attn_norm_result_golden[i*2048+j] - post_attn_norm_result[i*2048+j]);
                            if(post_attn_norm_result_golden[i*2048+j] != 0)
                                relative_error_temp =relative_error_temp + $abs(post_attn_norm_result_golden[i*2048+j] - post_attn_norm_result[i*2048+j]) / $abs(post_attn_norm_result_golden[i*2048+j]);
                        end
                        abs_error[i] = abs_error_temp/2048;
                        relative_error[i] = relative_error_temp/2048;
                        abs_error_temp = 0.0;
                        relative_error_temp = 0.0;
                    end
                    for (i =0 ; i< seq_len; i = i + 1) begin
                        $display("abs_error[%0d]: %f", i, abs_error[i]);
                        $display("relative_error[%0d]: %f", i, relative_error[i]);
                    end
                end
                default : begin
                    seq_len <= 7'd16;
                    post_attn_norm_hidden_size_cnt <= 1'b0;
                    start_post_attn_norm_residual <= 1'b0;
                    start_post_attn_norm_sqrt <= 1'b0;
                    post_attn_norm_ready <= 1'b0;
                    O_proj <= 1'b0;
                    Z0 <= 1'b0;
                    buffer_post_attn_norm_in <= 1'b0;
                    W_post_attn_norm <= 1'b0;
                    post_attn_norm_seq_cnt <= 1'b0;
                    state_select <= 1'b1;
                    post_attn_norm_decode_flag <= 1'b0;
                end
            endcase
        end
    end

    // ffn_residual fsm control
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            ffn_residual_ready <= 1'b0;
            start_ffn_residual <= 1'b0;
            D_proj             <= 1'b0;
            attn_residual_out  <= 1'b0;
            ffn_residual_hidden_size_cnt <= 1'b0;
        end 
        else begin
            case(state)
                IDLE: begin
                    ffn_residual_ready              <= 1'b0;
                    start_ffn_residual              <= 1'b0;
                    D_proj                          <= 1'b0;
                    attn_residual_out               <= 1'b0;
                    ffn_residual_hidden_size_cnt    <= 1'b0;
                end
                FFN_RESIDUAL : begin
                    if(!ffn_residual_ready) begin
                        start_ffn_residual <= 1'b1;
                        ffn_residual_ready <= 1'b1;
                        for(i = 0; i < M ; i = i + 1) begin
                            for(j = 0; j < N; j = j + 1) begin
                                D_proj[N*i*BW_FP + j*BW_FP +: BW_FP] <= down_proj[HIDDEN_SIZE*i + j + ffn_residual_hidden_size_cnt*N];
                                attn_residual_out[N*i*BW_FP + j*BW_FP +: BW_FP] <= attn_residual_result[HIDDEN_SIZE*i + j + ffn_residual_hidden_size_cnt*N];
                            end
                        end
                    end
                    else if(busy_ffn_residual_fall) begin
                        ffn_residual_ready <= 1'd0;
                        ffn_residual_hidden_size_cnt <= ffn_residual_hidden_size_cnt + 1'd1;
                    end
                    else begin
                        start_ffn_residual <= 1'b0;
                    end
                end
                FFN_RESIDUAL_CHECK: begin
                    for (i =0 ; i< 8; i = i + 1) begin
                        for(j = 0; j < 2048; j = j + 1) begin
                            $display("ffn_residual_result_golden[%0d]: %f", i*2048+j, ffn_residual_result_golden[i*2048+j]);
                            $display("ffn_residual_result[%0d]: %f", i*2048+j, ffn_residual_result[i*2048+j]);
                        end
                    end
                end
                default : begin
                    ffn_residual_ready              <= 1'b0;
                    start_ffn_residual              <= 1'b0;
                    D_proj                          <= 1'b0;
                    attn_residual_out               <= 1'b0;
                    ffn_residual_hidden_size_cnt    <= 1'b0;
                end
            endcase
        end
    end

    // ffn_mul fsm control
    always @(posedge clk or negedge rst_n) begin
        if(!rst_n) begin
            ffn_mul_ready <= 1'b0;
            start_ffn_mul <= 1'b0;
            U_proj        <= 1'b0;
            silu_in       <= 1'b0;
            ffn_mul_intermediate_size_cnt <= 1'b0;
        end 
        else begin
            case(state)
                IDLE: begin
                    ffn_mul_ready <= 1'b0;
                    start_ffn_mul <= 1'b0;
                    U_proj        <= 1'b0;
                    silu_in       <= 1'b0;
                    ffn_mul_intermediate_size_cnt <= 1'b0;
                end
                FFN_MUL : begin
                    if(!ffn_mul_ready) begin
                        start_ffn_mul <= 1'b1;
                        ffn_mul_ready <= 1'b1;
                        for(i = 0; i < M ; i = i + 1) begin
                            for(j = 0; j < N; j = j + 1) begin
                                U_proj[N*i*BW_FP + j*BW_FP +: BW_FP] <= up_proj[INTERMEDIATE_SIZE*i + j + ffn_mul_intermediate_size_cnt*N];
                                silu_in[N*i*BW_FP + j*BW_FP +: BW_FP] <= silu_gate[INTERMEDIATE_SIZE*i + j + ffn_mul_intermediate_size_cnt*N];
                            end
                        end
                    end
                    else if(busy_ffn_mul_fall) begin
                        ffn_mul_ready <= 1'd0;
                        ffn_mul_intermediate_size_cnt <= ffn_mul_intermediate_size_cnt + 1'd1;
                    end
                    else begin
                        start_ffn_mul <= 1'b0;
                    end
                end
                FFN_MUL_CHECK: begin
                    for (i =0 ; i< 8; i = i + 1) begin
                        for(j = 0; j < INTERMEDIATE_SIZE; j = j + 1) begin
                            $display("ffn_mul_golden[%0d]: %f", i*INTERMEDIATE_SIZE+j, ffn_mul_golden[i*INTERMEDIATE_SIZE+j]);
                            $display("ffn_mul_result[%0d]: %f", i*INTERMEDIATE_SIZE+j, ffn_mul_result[i*INTERMEDIATE_SIZE+j]);
                        end
                    end
                end
                default : begin
                    ffn_mul_ready <= 1'b0;
                    start_ffn_mul <= 1'b0;
                    U_proj        <= 1'b0;
                    silu_in       <= 1'b0;
                    ffn_mul_intermediate_size_cnt <= 1'b0;
                end
            endcase
        end
    end
/******************** test ****************************/ 
    // reg [16:0] dec_to_bf16_test;
    // real test_value_1;
    // real test_value_2;
    // real test_value_3;
    // initial begin
    //     dec_to_bf16_test = dec_to_bf16(5);
    //     $display("dec_to_bf16_test: %b", dec_to_bf16_test);
    //     test_value_1 = bf16_to_dec(17'h1f769);
    //     $display("test_value1: %f", test_value_1);
    //     test_value_2 = bf16_to_dec(17'h1f483);
    //     $display("test_value2: %f", test_value_2);
    //     test_value_3 = ffp_to_dec(29'hfe75500);
    //     $display("test_value3: %f", test_value_3);
    // end

/******************** initial ****************************/ 
	initial begin
		rst_n                   = 1'b0;
        rope_start              = 1'b0;
        post_attn_norm_start    = 1'b0;
        ffn_residual_start      = 1'b0;
        ffn_mul_start           = 1'b0;
		#(`clk_period*5 + 1);
        rst_n                   = 1'b1;
		#(`clk_period);
        rope_start              = 1'b0;
        post_attn_norm_start    = 1'b0;
        ffn_residual_start      = 1'b0;
        ffn_mul_start           = 1'b1;
        #(`clk_period);
        rope_start              = 1'b0;
        post_attn_norm_start    = 1'b0;
        ffn_residual_start      = 1'b0;
        ffn_mul_start           = 1'b0;
        #(`clk_period*20000);
		$finish;		
	end
	
    // clock generation
	initial clk= 1;
	always#(`clk_period/2) clk = ~clk;

    initial begin
        $fsdbDumpfile("tb_fma_top.fsdb");
        $fsdbDumpvars(0, tb_fma_top);
        $fsdbDumpMDA();
    end
    
/******************* BF16 convert function **********************************/
    function real two_pow;
        input integer e;    
        integer i;
        real r;
        begin
            r = 1.0;
            if (e >= 0) begin
                for (i = 0; i < e; i = i + 1) r = r * 2.0;
            end else begin
                for (i = 0; i < -e; i = i + 1) r = r / 2.0;
            end
            two_pow = r;
        end
    endfunction

    // Convert standard bfloat16 to decimal real number
    function real std_bf16_to_dec;
        input [15:0] bf; // 16-bit BF16 code
        // locals
        int    sign_bit;
        int    exp8;
        int    mant7;
        int    bias;
        real   sign;
        real   mant_frac;
        real   value;
        begin
            bias = 127; // bfloat16 uses bias 127
            sign_bit = bf[15];
            exp8 = bf[14:7];
            mant7 = bf[6:0];

            sign = (sign_bit == 1) ? -1.0 : 1.0;

            if (exp8 == 8'h00) begin
                // zero or subnormal
                if (mant7 == 0) begin
                    // +0 or -0
                    value = 0.0 * sign; // keep signed zero if simulator supports it
                end else begin
                    // subnormal: value = sign * 2^(1-bias) * (mant / 2^7)
                    mant_frac = (real'(mant7)) / (2.0 ** 7); // mant7/2^7
                    value = sign * two_pow(1 - bias) * mant_frac;
                end
            end else if (exp8 == 8'hFF) begin
                // infinity or NaN
                if (mant7 == 0) begin
                    // infinity
                    // 1.0/0.0 typically yields +Inf in simulators
                    value = sign * (1.0 / 0.0);
                end else begin
                    // NaN
                    value = 0.0 / 0.0; // yields NaN in most simulators
                end
            end else begin
                // normalized: value = sign * 2^(exp-bias) * (1 + mant/2^7)
                mant_frac = 1.0 + (real'(mant7)) / (2.0 ** 7);
                value = sign * two_pow(exp8 - bias) * mant_frac;
            end

            std_bf16_to_dec = value;
        end
    endfunction

    // Function to convert decimal value to BF16 format
    function [BW_FP-1:0] dec_to_bf16;  //{exp+2 ,comp {sign 1 m}}
        input real value;
        reg sign;
        integer exp_val;
        reg [7:0] exp_biased;
        reg [7:0] man_val;
        reg [8:0] man_twos;
        real abs_val, fraction;
        begin
            // Handle zero
            if (value == 0.0) begin
                dec_to_bf16 = {9'b0, 9'b0};
                return;
            end
            
            // Extract sign
            sign = (value < 0);
            abs_val = (value < 0) ? -value : value;
            
            // Calculate exponent
            exp_val = 0;
            if (abs_val >= 1.0) begin
                while (abs_val >= 2.0) begin
                    abs_val = abs_val / 2.0;
                    exp_val = exp_val + 1;
                end
            end else begin
                while (abs_val < 1.0) begin
                    abs_val = abs_val * 2.0;
                    exp_val = exp_val - 1;
                end
            end
            
            // Convert to biased exponent (subtract bias as requested)
            exp_biased = exp_val + 2;  // Note: subtracting bias as per your requirement
            
            // Calculate mantissa (fraction part)
            fraction = abs_val ;//- 1.0; // Remove the implicit 1
            man_val = $rtoi(fraction * 128.0); // Scale to 8-bit fraction
            
            // Convert to 9-bit two's complement
            if (sign) begin
                man_twos = ~{1'b0, man_val} + 1;
            end else begin
                man_twos = {1'b0, man_val};
            end
            
            // Pack into BF16 format: [17:9] = exponent, [8:0] = mantissa
            dec_to_bf16 = {exp_biased, man_twos};
        end
    endfunction


  function real bf16_to_dec;
      input [BW_FP - 1:0] bf16_val;
      reg sign;
      real exp_val,exp_abs;
      reg [7:0] man_val;
      real fraction, result;
      begin
          // Extract components
          if (bf16_val[16]) begin
              // Negative: convert from two's complement
              exp_abs = $itor((~bf16_val[16:9] + 1) & 8'hFF) ;
              exp_val = -exp_abs ;
          end else begin
              // Positive
              exp_abs = $itor(bf16_val[16:9]) ;
              exp_val = exp_abs ;
          end
          //exp_val = $signed(bf16_val[16:9]);// + BIAS; // Add back bias
        
          man_val = bf16_val[7:0];
          sign = bf16_val[8]; // Sign bit is MSB of mantissa field
          
          // Handle zero
          if (bf16_val == 0) begin
              bf16_to_dec = 0.0;
              return;
          end
  
          if (sign) begin
              // Negative: convert from two's complement
              fraction = $itor((~{sign, man_val} + 1) & 9'h1FF) / 512.0;
          end else begin
              // Positive
              fraction = $itor(man_val) / 512.0;
          end

          result = (/*1.0 +*/ fraction) * (2.0 ** exp_val);
          bf16_to_dec = sign ? -result : result;
      end
  endfunction


  function real ffp_to_dec;
      input [28:0] bf16_val;
      reg sign;
      real exp_val,exp_abs;
      reg [17:0] man_val;
      real fraction, result;
      begin
          // Extract components
          if (bf16_val[28]) begin
              // Negative: convert from two's complement
              exp_abs = $itor((~bf16_val[28:19] + 1) & 10'h1FF) ;
              exp_val = -exp_abs ;
          end else begin
              // Positive
              exp_abs = $itor(bf16_val[28:19]) ;
              exp_val = exp_abs ;
          end
                  
          man_val = bf16_val[17:0];
          sign = bf16_val[18]; 

          // Handle zero
          if (bf16_val == 0) begin
              ffp_to_dec = 0.0;
              return;
          end
  
          if (sign) begin
              // Negative: convert from two's complement
              fraction = $itor((~{sign, man_val} + 1) & 19'h7FFFF) / (2**19);
          end else begin
              // Positive
              fraction = $itor(man_val) / (2**19);
          end

          result = (/*1.0 +*/ fraction) * (2.0 ** exp_val);
          ffp_to_dec = sign ? -result : result;
      end
  endfunction
endmodule
